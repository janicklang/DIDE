library ieee;
use ieee.std_logic_1164.all;

entity MyAnd is

end MyAnd;

architecture rtl of MyAnd is
  
begin
  
end rtl;
