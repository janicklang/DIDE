library ieee;
use ieee.std_logic_1164.all;

entity MyNand is
  port(
    u_pi : in  std_logic;
    v_pi : in  std_logic;
    w_po : out std_logic
    );
end MyNand;

architecture struct of MyNand is

begin

end struct;
