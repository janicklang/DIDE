library ieee;
use ieee.std_logic_1164.all;

entity MyInv is

end MyInv;

architecture rtl of MyInv is
  
begin
  
end rtl;
